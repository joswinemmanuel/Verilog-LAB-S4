`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:17:30 06/09/2023 
// Design Name: 
// Module Name:    Logic_gates_structural 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module Logic_gates_structural(
    input a,
    input b,
    output c_and,
    output c_or,
    output c_not,
    output c_xor,
    output c_nand,
    output c_nor,
    output c_xnor
    );
  
	 and(c_and, a, b);
	 or(c_or, a, b);
	 not(c_not, a, b);
	 xor(c_xor, a, b);
	 nand(c_nand, a, b);
	 nor(c_nor, a, b);
	 xnor(c_xnor, a, b);
  
endmodule
